`include "head.v"



